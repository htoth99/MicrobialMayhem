system.number,seqid,system,target.name,hmm.accession,hmm.name,protein.name,full.seq.E.value,domain.iE.value,target.coverage,hmm.coverage,start,end,strand,target.description,relative.position,contig.end,all.domains,best.hits
1,NZ_CP025084.1,cas_type_I-E,WP_037380268.1,PDLC01768,Cas3e_WP_058658455.1,Cas3e,7.499999999999996e-215,7.499999999999996e-215,0.603,0.991,1077064,1079808,+,CRISPR-associated helicase/endonuclease Cas3 [Serratia sp. ATCC 39006],960,4398,"PDLC01767,Cas3e_WP_189128522.1, 1, 1.2e-213, 0.979, 0.921 | PDLC01768,Cas3e_WP_058658455.1, 1, 190, 0.05, 0.083 | PDLC01768,Cas3e_WP_058658455.1, 2, 7.5e-215, 0.603, 0.991","PDLC01768, Cas3e_WP_058658455.1, 7.5e-215, 0.603, 0.991 | PDLC01767, Cas3e_WP_189128522.1, 1.2e-213, 0.979, 0.921"
1,NZ_CP025084.1,cas_type_I-E,WP_021013291.1,PDLC00999,casA_cse1,Cas8e,3.599999999999999e-135,4.299999999999999e-135,0.959,0.994,1079875,1081416,+,type I-E CRISPR-associated protein Cse1/CasA [Serratia sp. ATCC 39006],961,4398,"PDLC00999,casA_cse1, 1, 4.3e-135, 0.959, 0.994 | PDLC01282,cd09669, 1, 5.9e-125, 0.957, 0.993 | PDLC01342,cd09729, 1, 5e-118, 0.901, 0.998 | PDLC01622,pfam09481, 1, 2.3e-105, 0.869, 0.986","PDLC00999, casA_cse1, 4.3e-135, 0.959, 0.994 | PDLC01282, cd09669, 5.9e-125, 0.957, 0.993 | PDLC01342, cd09729, 5e-118, 0.901, 0.998 | PDLC01622, pfam09481, 2.3e-105, 0.869, 0.986"
1,NZ_CP025084.1,cas_type_I-E,WP_021013290.1,PDLC01000,casB_cse2,Cas11e,1.7e-28,1.9e-28,0.807,0.962,1081409,1082032,+,type I-E CRISPR-associated protein Cse2/CasB [Serratia sp. ATCC 39006],962,4398,"PDLC01000,casB_cse2, 1, 1.9e-28, 0.807, 0.962 | PDLC01283,cd09670, 1, 8.2e-25, 0.792, 0.929 | PDLC01344,cd09731, 1, 2.1e-23, 0.729, 0.977 | PDLC01624,pfam09485, 1, 3e-18, 0.72, 0.984","PDLC01000, casB_cse2, 1.9e-28, 0.807, 0.962 | PDLC01283, cd09670, 8.2e-25, 0.792, 0.929 | PDLC01344, cd09731, 2.1e-23, 0.729, 0.977 | PDLC01624, pfam09485, 3e-18, 0.72, 0.984"
1,NZ_CP025084.1,cas_type_I-E,WP_021013289.1,PDLC00959,casC_Cse4,Cas7e,1.5999999999999996e-101,1.7999999999999997e-101,0.912,0.997,1082035,1083093,+,type I-E CRISPR-associated protein Cas7/Cse4/CasC [Serratia sp. ATCC 39006],963,4398,"PDLC00959,casC_Cse4, 1, 1.8e-101, 0.912, 0.997 | PDLC01259,cd09646, 1, 6.5e-95, 0.912, 0.997 | PDLC01620,pfam09344, 1, 4.6e-96, 0.952, 0.955","PDLC00959, casC_Cse4, 1.8e-101, 0.912, 0.997 | PDLC01620, pfam09344, 4.6e-96, 0.952, 0.955 | PDLC01259, cd09646, 6.5e-95, 0.912, 0.997"
1,NZ_CP025084.1,cas_type_I-E,WP_021013288.1,PDLC00949,casD_Cas5e,Cas5e,2.8999999999999998e-52,3.2999999999999996e-52,0.947,0.978,1083105,1083839,+,type I-E CRISPR-associated protein Cas5/CasD [Serratia sp. ATCC 39006],964,4398,"PDLC00949,casD_Cas5e, 1, 3.3e-52, 0.947, 0.978 | PDLC01258,cd09645, 1, 2.4e-50, 0.672, 0.873 | PDLC01369,cd09756, 1, 3.6e-49, 0.672, 0.871","PDLC00949, casD_Cas5e, 3.3e-52, 0.947, 0.978 | PDLC01258, cd09645, 2.4e-50, 0.672, 0.873 | PDLC01369, cd09756, 3.6e-49, 0.672, 0.871"
1,NZ_CP025084.1,cas_type_I-E,WP_021013287.1,PDLC00954,casE_Cse3,Cas6e,7.399999999999999e-60,8.2e-60,0.991,0.99,1083839,1084486,+,type I-E CRISPR-associated protein Cas6/Cse3/CasE [Serratia sp. ATCC 39006],965,4398,"PDLC00954,casE_Cse3, 1, 8.2e-60, 0.991, 0.99 | PDLC01277,cd09664, 1, 4.9e-54, 0.967, 0.994 | PDLC01340,cd09727, 1, 3.1e-51, 0.991, 0.995","PDLC00954, casE_Cse3, 8.2e-60, 0.991, 0.99 | PDLC01277, cd09664, 4.9e-54, 0.967, 0.994 | PDLC01340, cd09727, 3.1e-51, 0.991, 0.995"
1,NZ_CP025084.1,cas_type_I-E,WP_021013286.1,PDLC01744,Cas1e_WP_035839043.1,Cas1e,3.499999999999999e-118,3.999999999999999e-118,0.879,0.866,1084510,1085433,+,type I-E CRISPR-associated endonuclease Cas1e [Serratia sp. ATCC 39006],966,4398,"PDLC00924,cas1_ECOLI, 1, 3.6e-114, 0.86, 0.985 | PDLC01744,Cas1e_WP_035839043.1, 1, 4e-118, 0.879, 0.866 | PDLC01745,Cas1e_WP_120372217.1, 1, 1.2e-63, 0.86, 0.941 | PDLC01746,Cas1e_WP_162621937.1, 1, 3.5e-81, 0.524, 0.994","PDLC01744, Cas1e_WP_035839043.1, 4e-118, 0.879, 0.866 | PDLC00924, cas1_ECOLI, 3.6e-114, 0.86, 0.985 | PDLC01746, Cas1e_WP_162621937.1, 3.5e-81, 0.524, 0.994 | PDLC01745, Cas1e_WP_120372217.1, 1.2e-63, 0.86, 0.941"
1,NZ_CP025084.1,cas_type_I-E,WP_021013285.1,PDLC01752,Cas2e_WP_051024046.1,Cas2e,1.9e-44,2.1e-44,0.938,0.783,1085430,1085723,+,type I-E CRISPR-associated endoribonuclease Cas2 [Serratia sp. ATCC 39006],967,4398,"PDLC00934,cas_CT1978, 1, 1.3e-40, 0.876, 0.989 | PDLC01752,Cas2e_WP_051024046.1, 1, 2.1e-44, 0.938, 0.783 | PDLC01753,Cas2e_WP_128219160.1, 1, 1.2e-28, 0.938, 0.892 | PDLC01754,Cas2e_WP_012568472.1, 1, 2.6e-16, 0.907, 0.959 | PDLC01755,Cas2e_WP_081586257.1, 1, 1.5e-13, 0.897, 0.632","PDLC01752, Cas2e_WP_051024046.1, 2.1e-44, 0.938, 0.783 | PDLC00934, cas_CT1978, 1.3e-40, 0.876, 0.989 | PDLC01753, Cas2e_WP_128219160.1, 1.2e-28, 0.938, 0.892 | PDLC01754, Cas2e_WP_012568472.1, 2.6e-16, 0.907, 0.959 | PDLC01755, Cas2e_WP_081586257.1, 1.5e-13, 0.897, 0.632"
4,NZ_CP025084.1,CRISPR_array,CRISPR001,NA,NA,CRISPR_array,NA,6.25,NA,NA,1085808,1089009,+,CRISPR001; repeat=GTGTTCCCCGCACCCGCGGGGATAAACCG; score=6.25,967.01,4398,NA,NA
2,NZ_CP025084.1,cas_type_I-F1,WP_021017054.1,PDLC01352,cd09739,Cas6f,1.0999999999999999e-67,1.3e-67,0.995,0.995,1426973,1427527,-,type I-F CRISPR-associated endoribonuclease Cas6/Csy4 [Serratia sp. ATCC 39006],1255,4398,"PDLC00955,cas_Csy4, 1, 6.4e-57, 0.984, 0.995 | PDLC01287,cd09674, 1, 1.5e-61, 0.995, 0.995 | PDLC01352,cd09739, 1, 1.3e-67, 0.995, 0.995 | PDLC01631,pfam09618, 1, 7.1e-66, 0.978, 0.994","PDLC01352, cd09739, 1.3e-67, 0.995, 0.995 | PDLC01631, pfam09618, 7.1e-66, 0.978, 0.994 | PDLC01287, cd09674, 1.5e-61, 0.995, 0.995 | PDLC00955, cas_Csy4, 6.4e-57, 0.984, 0.995"
2,NZ_CP025084.1,cas_type_I-F1,WP_021017053.1,PDLC01629,pfam09615,Cas7f,3.299999999999999e-146,3.699999999999999e-146,0.961,0.997,1427537,1428544,-,type I-F CRISPR-associated protein Csy3 [Serratia sp. ATCC 39006],1256,4398,"PDLC01030,cas_Csy3, 1, 3.2e-140, 0.973, 0.997 | PDLC01290,cd09677, 1, 2e-135, 0.973, 0.997 | PDLC01350,cd09737, 1, 3.7e-140, 0.964, 0.997 | PDLC01629,pfam09615, 1, 3.7e-146, 0.961, 0.997","PDLC01629, pfam09615, 3.7e-146, 0.961, 0.997 | PDLC01030, cas_Csy3, 3.2e-140, 0.973, 0.997 | PDLC01350, cd09737, 3.7e-140, 0.964, 0.997 | PDLC01290, cd09677, 2e-135, 0.973, 0.997"
2,NZ_CP025084.1,cas_type_I-F1,WP_021017052.1,PDLC01029,cas_Csy2,Cas5f,7.299999999999998e-118,8.299999999999998e-118,0.926,0.993,1428555,1429490,-,type I-F CRISPR-associated protein Csy2 [Serratia sp. ATCC 39006],1257,4398,"PDLC01029,cas_Csy2, 1, 8.3e-118, 0.926, 0.993 | PDLC01199,C19_Cas5f_1, 1, 2e-07, 0.418, 0.506 | PDLC01199,C19_Cas5f_1, 2, 0.054, 0.196, 0.232 | PDLC01289,cd09676, 1, 2.8e-110, 0.926, 0.992 | PDLC01349,cd09736, 1, 4.8e-92, 0.923, 0.992 | PDLC01628,pfam09614, 1, 1.4e-99, 0.923, 0.996","PDLC01029, cas_Csy2, 8.3e-118, 0.926, 0.993 | PDLC01289, cd09676, 2.8e-110, 0.926, 0.992 | PDLC01628, pfam09614, 1.4e-99, 0.923, 0.996 | PDLC01349, cd09736, 4.8e-92, 0.923, 0.992 | PDLC01199, C19_Cas5f_1, 2e-07, 0.418, 0.506"
2,NZ_CP025084.1,cas_type_I-F1,WP_021017051.1,PDLC01028,cas_Csy1,Cas8f,3.299999999999999e-158,3.999999999999999e-158,0.847,0.997,1429487,1430821,-,type I-F CRISPR-associated protein Csy1 [Serratia sp. ATCC 39006],1258,4398,"PDLC01028,cas_Csy1, 1, 4e-158, 0.847, 0.997 | PDLC01288,cd09675, 1, 9.5e-152, 0.847, 0.997 | PDLC01348,cd09735, 1, 7.6e-140, 0.822, 0.994 | PDLC01627,pfam09611, 1, 3.2e-133, 0.82, 0.994","PDLC01028, cas_Csy1, 4e-158, 0.847, 0.997 | PDLC01288, cd09675, 9.5e-152, 0.847, 0.997 | PDLC01348, cd09735, 7.6e-140, 0.822, 0.994 | PDLC01627, pfam09611, 3.2e-133, 0.82, 0.994"
2,NZ_CP025084.1,cas_type_I-F1,WP_021017050.1,PDLC00941,cas3_yersinia,Cas23f,0,0,0.997,0.999,1430845,1434129,-,type I-F CRISPR-associated helicase Cas3f [Serratia sp. ATCC 39006],1259,4398,"PDLC00941,cas3_yersinia, 1, 0, 0.997, 0.999","PDLC00941, cas3_yersinia, 0, 0.997, 0.999"
2,NZ_CP025084.1,cas_type_I-F1,WP_021017049.1,PDLC00925,cas1_YPEST,Cas1f,4.399999999999998e-159,5.099999999999997e-159,0.936,0.993,1434126,1435106,-,type I-F CRISPR-associated endonuclease Cas1f [Serratia sp. ATCC 39006],1260,4398,"PDLC00925,cas1_YPEST, 1, 5.1e-159, 0.936, 0.993","PDLC00925, cas1_YPEST, 5.1e-159, 0.936, 0.993"
4,NZ_CP025084.1,CRISPR_array,CRISPR002,NA,NA,CRISPR_array,NA,6.24,NA,NA,1435404,1438854,+,CRISPR002; repeat=GTTCACTGCCGTACAGGCAGCTTAGAAA; score=6.24,1260.02,4398,NA,NA
3,NZ_CP025084.1,cas_type_III-A,WP_021014796.1,PDLC01248,cd09634,Cas1,1.5e-44,1.7e-44,0.969,0.976,4374503,4375384,+,CRISPR-associated endonuclease Cas1 [Serratia sp. ATCC 39006],3843,4398,"PDLC00922,cas1_MYXAN, 1, 0.037, 0.338, 0.288 | PDLC00922,cas1_MYXAN, 2, 2e-09, 0.297, 0.265 | PDLC00923,cas1_DVULG, 1, 1.1e-08, 0.399, 0.35 | PDLC00923,cas1_DVULG, 2, 3e-15, 0.423, 0.382 | PDLC00924,cas1_ECOLI, 1, 0.00018, 0.321, 0.357 | PDLC00924,cas1_ECOLI, 2, 9.6, 0.184, 0.193 | PDLC00926,cas1_NMENI, 1, 4.3e-13, 0.785, 0.827 | PDLC00927,cas1, 1, 9.6e-35, 0.904, 0.881 | PDLC00928,cas1_I_II_III_V_maka, 1, 4e-34, 0.976, 0.984 | PDLC00929,cas1_PREFRAN, 1, 16, 0.273, 0.246 | PDLC00929,cas1_PREFRAN, 2, 5.4e-10, 0.478, 0.432 | PDLC01248,cd09634, 1, 1.7e-44, 0.969, 0.976 | PDLC01249,cd09636, 1, 8.1e-32, 0.809, 0.988 | PDLC01332,cd09719, 1, 0.00036, 0.321, 0.364 | PDLC01332,cd09719, 2, 8.7, 0.184, 0.199 | PDLC01333,cd09720, 1, 8.1e-14, 0.775, 0.833 | PDLC01334,cd09721, 1, 5.8e-08, 0.403, 0.354 | PDLC01334,cd09721, 2, 1.7e-15, 0.423, 0.387 | PDLC01335,cd09722, 1, 2.4e-21, 0.816, 0.794 | PDLC01449,COG1518, 1, 4.6e-35, 0.98, 0.947 | PDLC01608,pfam01867, 1, 2.1e-41, 0.881, 0.982 | PDLC01740,Cas1_IIIa_WP_158094482.1, 1, 300, 0.184, 0.157 | PDLC01740,Cas1_IIIa_WP_158094482.1, 2, 1.8e-12, 0.416, 0.378 | PDLC01741,Cas1_IIIa_WP_000655858.1, 1, 0.019, 0.727, 0.711 | PDLC01742,Cas1b_WP_142933338.1, 1, 1.4e-23, 0.863, 0.822 | PDLC01743,Cas1c_WP_008519397.1, 1, 3.8e-08, 0.406, 0.356 | PDLC01743,Cas1c_WP_008519397.1, 2, 4.7e-18, 0.427, 0.386 | PDLC01744,Cas1e_WP_035839043.1, 1, 0.0093, 0.283, 0.278 | PDLC01744,Cas1e_WP_035839043.1, 2, 100, 0.184, 0.17 | PDLC01745,Cas1e_WP_120372217.1, 1, 0.0023, 0.3, 0.319 | PDLC01745,Cas1e_WP_120372217.1, 2, 220, 0.085, 0.08 | PDLC01747,Cas1g_WP_005511840.1, 1, 3.8e-20, 0.853, 0.509 | PDLC02025,Cas1d_Cas1d, 1, 6.3e-28, 0.898, 0.851 | PDLC02061,Cas1_II_WP_078484493.1, 1, 1.6e-14, 0.805, 0.657 | PDLC02062,Cas1_II_WP_122951193.1, 1, 0.00024, 0.369, 0.344 | PDLC02062,Cas1_II_WP_122951193.1, 2, 1.8e-05, 0.311, 0.29 | PDLC02062,Cas1_II_WP_122951193.1, 3, 500, 0.048, 0.044 | PDLC02063,Cas1_IIIb_Cas1_IIIb, 1, 7.6e-14, 0.809, 0.397 | PDLC02064,Cas1a_Cas1a, 1, 1.2e-09, 0.785, 0.816 | PDLC02065,Cas1b_WP_013704840.1, 1, 3.4e-19, 0.457, 0.41 | PDLC02066,Cas1b_WP_035727688.1, 1, 0.042, 0.396, 0.363 | PDLC02066,Cas1b_WP_035727688.1, 2, 5.2e-14, 0.553, 0.5 | PDLC02067,Cas1b_WP_188882336.1, 1, 0.005, 0.355, 0.197 | PDLC02067,Cas1b_WP_188882336.1, 2, 4e-10, 0.406, 0.233","PDLC01248, cd09634, 1.7e-44, 0.969, 0.976 | PDLC01608, pfam01867, 2.1e-41, 0.881, 0.982 | PDLC01449, COG1518, 4.6e-35, 0.98, 0.947 | PDLC00927, cas1, 9.6e-35, 0.904, 0.881 | PDLC00928, cas1_I_II_III_V_maka, 4e-34, 0.976, 0.984"
3,NZ_CP025084.1,cas_type_III-A,WP_021014795.1,PDLC01338,cd09725,Cas2,8e-12,9.9e-12,0.663,0.816,4375377,4375673,+,CRISPR-associated endonuclease Cas2 [Serratia sp. ATCC 39006],3844,4398,"PDLC00935,cas2, 1, 4.4e-07, 0.653, 0.708 | PDLC00936,cas2_I_II_III_V_maka, 1, 9e-08, 0.633, 0.783 | PDLC01251,cd09638, 1, 9.4e-07, 0.643, 0.738 | PDLC01338,cd09725, 1, 9.9e-12, 0.663, 0.816 | PDLC01443,COG1343, 1, 1.1e-07, 0.663, 0.733 | PDLC01525,mkCas0128, 1, 0.014, 0.622, 0.678 | PDLC01649,pfam09827, 1, 3.6e-09, 0.653, 0.9 | PDLC01748,Cas2_IIIa_Cas2_IIIa, 1, 9.8e-06, 0.592, 0.648 | PDLC01749,Cas2b_WP_014295803.1, 1, 0.00017, 0.612, 0.678 | PDLC01751,Cas2c_WP_035173219.1, 1, 4.8e-07, 0.571, 0.642 | PDLC01756,Cas2g_WP_109723797.1, 1, 1.9e-10, 0.663, 0.677 | PDLC02027,Cas2d_WP_013277804.1, 1, 7.1e-06, 0.622, 0.685 | PDLC02070,Cas2_II_WP_021888968.1, 1, 4.4e-05, 0.643, 0.708 | PDLC02074,Cas2_IIIb_Cas2_IIIb, 1, 5.2e-06, 0.633, 0.709 | PDLC02076,Cas2b_WP_066217071.1, 1, 0.0051, 0.582, 0.644 | PDLC02077,Cas2b_WP_028460064.1, 1, 5.7e-06, 0.663, 0.677 | PDLC02078,Cas2b_WP_038071942.1, 1, 9.9e-11, 0.673, 0.691","PDLC01338, cd09725, 9.9e-12, 0.663, 0.816 | PDLC02078, Cas2b_WP_038071942.1, 9.9e-11, 0.673, 0.691 | PDLC01756, Cas2g_WP_109723797.1, 1.9e-10, 0.663, 0.677 | PDLC01649, pfam09827, 3.6e-09, 0.653, 0.9 | PDLC00936, cas2_I_II_III_V_maka, 9e-08, 0.633, 0.783"
4,NZ_CP025084.1,CRISPR_array,CRISPR003,NA,NA,CRISPR_array,NA,6.08,NA,NA,4375925,4376651,+,CRISPR003; repeat=GTCCTTACGGACGCTCCCTGACTGAAGGGATTAAGAC; score=6.08,3844.03,4398,NA,NA
3,NZ_CP025084.1,cas_type_III-A,WP_021014794.1,PDLC00916,cas_TM1811_Csm1,Cas10a,4.999999999999999e-90,1.1999999999999997e-89,0.681,0.783,4376785,4379235,+,type III-A CRISPR-associated protein Cas10/Csm1 [Serratia sp. ATCC 39006],3845,4398,"PDLC00916,cas_TM1811_Csm1, 1, 1.2e-89, 0.681, 0.783 | PDLC00916,cas_TM1811_Csm1, 2, 840, 0.059, 0.068 | PDLC00919,cas10_III_maka_5, 1, 14, 0.168, 0.312 | PDLC00919,cas10_III_maka_5, 2, 2.1e-05, 0.083, 0.184 | PDLC01292,cd09679, 1, 2.4e-07, 0.168, 0.326 | PDLC01293,cd09680, 1, 4.2e-87, 0.691, 0.808 | PDLC01422,cls000742, 1, 2.2e-07, 0.261, 0.401 | PDLC01444,COG1353, 1, 2e-16, 0.344, 0.336 | PDLC01444,COG1353, 2, 6.6e-26, 0.272, 0.336 | PDLC01529,mkCas0133, 1, 28, 0.165, 0.314 | PDLC01529,mkCas0133, 2, 3.7e-06, 0.086, 0.192 | PDLC01739,Cas10_IIIa_WP_087192840.1, 1, 3.1e-19, 0.283, 0.317 | PDLC01739,Cas10_IIIa_WP_087192840.1, 2, 3.4e-26, 0.32, 0.319","PDLC00916, cas_TM1811_Csm1, 1.2e-89, 0.681, 0.783 | PDLC01293, cd09680, 4.2e-87, 0.691, 0.808 | PDLC01739, Cas10_IIIa_WP_087192840.1, 3.4e-26, 0.32, 0.319 | PDLC01444, COG1353, 6.6e-26, 0.272, 0.336 | PDLC01422, cls000742, 2.2e-07, 0.261, 0.401"
3,NZ_CP025084.1,cas_type_III-A,WP_021014793.1,PDLC01612,pfam03750,Csm2,9.4e-16,1.2e-15,0.78,0.921,4379260,4379643,+,type III-A CRISPR-associated protein Csm2 [Serratia sp. ATCC 39006],3846,4398,"PDLC01010,cas_TM1810_Csm2, 1, 2600, 0, 0 | PDLC01010,cas_TM1810_Csm2, 2, 1.5e-14, 0.685, 0.969 | PDLC01012,csm2_IIIA_maka_7, 1, 1.7e-07, 0.717, 0.662 | PDLC01260,cd09647, 1, 2.5e-14, 0.677, 0.965 | PDLC01433,cls001490, 1, 0.005, 0.276, 0.182 | PDLC01446,COG1421, 1, 3.8e-11, 0.921, 0.785 | PDLC01547,mkCas0157, 1, 0.0013, 0.732, 0.74 | PDLC01576,mkCas0187, 1, 7.4e-07, 0.661, 0.874 | PDLC01612,pfam03750, 1, 1.2e-15, 0.78, 0.921","PDLC01612, pfam03750, 1.2e-15, 0.78, 0.921 | PDLC01010, cas_TM1810_Csm2, 1.5e-14, 0.685, 0.969 | PDLC01260, cd09647, 2.5e-14, 0.677, 0.965 | PDLC01446, COG1421, 3.8e-11, 0.921, 0.785 | PDLC01012, csm2_IIIA_maka_7, 1.7e-07, 0.717, 0.662"
3,NZ_CP025084.1,cas_type_III-A,WP_021014792.1,PDLC01297,cd09684,Csm3,9.4e-61,1.3e-60,0.887,0.955,4379656,4380402,+,type III-A CRISPR-associated RAMP protein Csm3 [Serratia sp. ATCC 39006],3847,4398,"PDLC00981,cas_RAMP_Cmr4, 1, 1.2e-09, 0.202, 0.17 | PDLC00981,cas_RAMP_Cmr4, 2, 190, 0.077, 0.067 | PDLC00982,cmr4_IIIB_maka, 1, 5.1e-09, 0.202, 0.171 | PDLC00982,cmr4_IIIB_maka, 2, 960, 0.065, 0.057 | PDLC01013,csm3_IIIAD_maka_1, 1, 0.00059, 0.202, 0.077 | PDLC01014,cas7_TM1809, 1, 2.4e-60, 0.855, 0.975 | PDLC01015,csm3_IIID_maka_5, 1, 1.8e-10, 0.802, 0.983 | PDLC01016,csm3_IIIAD_maka_5, 1, 1.1e-10, 0.835, 0.989 | PDLC01017,csm3_IIID_maka_6, 1, 8.2e-44, 0.875, 0.817 | PDLC01018,cas5_csm4, 1, 0.012, 0.129, 0.106 | PDLC01019,csm4_IIIA_maka_3, 1, 0.0098, 0.145, 0.119 | PDLC01020,cas_TM1807_csm5, 1, 0.00011, 0.085, 0.058 | PDLC01021,csm5_IIIA_maka_3, 1, 1000, 0.056, 0.038 | PDLC01021,csm5_IIIA_maka_3, 2, 0.00055, 0.109, 0.07 | PDLC01024,cas_cyan_RAMP_2, 1, 19, 0.081, 0.05 | PDLC01024,cas_cyan_RAMP_2, 2, 0.018, 0.157, 0.095 | PDLC01130,icity0028, 1, 290, 0.109, 0.092 | PDLC01130,icity0028, 2, 0.015, 0.286, 0.224 | PDLC01275,cd09662, 1, 2.7e-05, 0.109, 0.078 | PDLC01276,cd09663, 1, 940, 0.085, 0.078 | PDLC01276,cd09663, 2, 0.009, 0.117, 0.108 | PDLC01295,cd09682, 1, 2.1e-09, 0.218, 0.176 | PDLC01295,cd09682, 2, 110, 0.21, 0.195 | PDLC01296,cd09683, 1, 1.5e-11, 0.867, 0.958 | PDLC01297,cd09684, 1, 1.3e-60, 0.887, 0.955 | PDLC01313,cd09700, 1, 15, 0.089, 0.065 | PDLC01313,cd09700, 2, 0.07, 0.153, 0.086 | PDLC01339,cd09726, 1, 2.1e-09, 0.218, 0.258 | PDLC01339,cd09726, 2, 2400, 0.089, 0.129 | PDLC01339,cd09726, 3, 0.077, 0.222, 0.27 | PDLC01407,cls000253, 1, 0.00013, 0.21, 0.092 | PDLC01407,cls000253, 2, 28, 0.282, 0.131 | PDLC01420,cls000715, 1, 24, 0.077, 0.055 | PDLC01420,cls000715, 2, 0.04, 0.129, 0.082 | PDLC01440,Csm5, 1, 230, 0.06, 0.047 | PDLC01440,Csm5, 2, 1.7e-05, 0.117, 0.084 | PDLC01441,COG1336, 1, 3.8e-09, 0.198, 0.184 | PDLC01441,COG1336, 2, 100, 0.218, 0.204 | PDLC01442,COG1337, 1, 1e-43, 0.903, 0.88 | PDLC01450,COG1567, 1, 0.0018, 0.153, 0.141 | PDLC01571,mkCas0182, 1, 980, 0.069, 0.05 | PDLC01571,mkCas0182, 2, 0.01, 0.069, 0.05 | PDLC01585,mkCas0198, 1, 0.51, 0.194, 0.218 | PDLC01585,mkCas0198, 2, 13, 0.133, 0.16 | PDLC01613,pfam03787, 1, 1e-11, 0.835, 0.994 | PDLC01733,COG1332, 1, 1100, 0.056, 0.038 | PDLC01733,COG1332, 2, 8.3e-06, 0.113, 0.07","PDLC01297, cd09684, 1.3e-60, 0.887, 0.955 | PDLC01014, cas7_TM1809, 2.4e-60, 0.855, 0.975 | PDLC01017, csm3_IIID_maka_6, 8.2e-44, 0.875, 0.817 | PDLC01442, COG1337, 1e-43, 0.903, 0.88 | PDLC01613, pfam03787, 1e-11, 0.835, 0.994"
3,NZ_CP025084.1,cas_type_III-A,WP_021014791.1,PDLC01494,mkCas0089,Csm4,2.0999999999999999e-97,2.4e-97,0.945,0.99,4380402,4381382,+,hypothetical protein [Serratia sp. ATCC 39006],3848,4398,"PDLC01018,cas5_csm4, 1, 0.0079, 0.245, 0.258 | PDLC01276,cd09663, 1, 4.9e-08, 0.693, 0.78 | PDLC01450,COG1567, 1, 3.4e-05, 0.641, 0.73 | PDLC01494,mkCas0089, 1, 2.4e-97, 0.945, 0.99","PDLC01494, mkCas0089, 2.4e-97, 0.945, 0.99 | PDLC01276, cd09663, 4.9e-08, 0.693, 0.78 | PDLC01450, COG1567, 3.4e-05, 0.641, 0.73 | PDLC01018, cas5_csm4, 0.0079, 0.245, 0.258"
3,NZ_CP025084.1,cas_type_III-A,WP_021014790.1,PDLC01440,Csm5,Csm5,5.1e-18,1.3e-17,0.705,0.981,4381379,4383058,+,DUF324 domain-containing protein [Serratia sp. ATCC 39006],3849,4398,"PDLC00916,cas_TM1811_Csm1, 1, 0.036, 0.17, 0.145 | PDLC00981,cas_RAMP_Cmr4, 1, 75, 0.029, 0.057 | PDLC00981,cas_RAMP_Cmr4, 2, 0.0062, 0.055, 0.095 | PDLC00981,cas_RAMP_Cmr4, 3, 920, 0.077, 0.159 | PDLC00982,cmr4_IIIB_maka, 1, 27, 0.03, 0.06 | PDLC00982,cmr4_IIIB_maka, 2, 0.0036, 0.052, 0.089 | PDLC01013,csm3_IIIAD_maka_1, 1, 0.05, 0.034, 0.029 | PDLC01014,cas7_TM1809, 1, 0.0026, 0.063, 0.172 | PDLC01015,csm3_IIID_maka_5, 1, 3900, 0.023, 0.073 | PDLC01015,csm3_IIID_maka_5, 2, 0.00084, 0.039, 0.107 | PDLC01016,csm3_IIIAD_maka_5, 1, 1.6e-05, 0.277, 0.307 | PDLC01017,csm3_IIID_maka_6, 1, 2.4e-05, 0.045, 0.097 | PDLC01020,cas_TM1807_csm5, 1, 6.6, 0.045, 0.069 | PDLC01020,cas_TM1807_csm5, 2, 6.5e-10, 0.175, 0.258 | PDLC01020,cas_TM1807_csm5, 3, 2300, 0.048, 0.077 | PDLC01021,csm5_IIIA_maka_3, 1, 150, 0.043, 0.064 | PDLC01021,csm5_IIIA_maka_3, 2, 1.4e-07, 0.165, 0.239 | PDLC01021,csm5_IIIA_maka_3, 3, 1700, 0.038, 0.056 | PDLC01275,cd09662, 1, 2.5e-12, 0.358, 0.52 | PDLC01275,cd09662, 2, 1100, 0.055, 0.087 | PDLC01295,cd09682, 1, 110, 0.03, 0.066 | PDLC01295,cd09682, 2, 0.017, 0.047, 0.102 | PDLC01296,cd09683, 1, 0.01, 0.064, 0.203 | PDLC01297,cd09684, 1, 0.0039, 0.048, 0.126 | PDLC01339,cd09726, 1, 7.8e-06, 0.1, 0.294 | PDLC01407,cls000253, 1, 0.0039, 0.054, 0.058 | PDLC01407,cls000253, 2, 980, 0.032, 0.035 | PDLC01440,Csm5, 1, 1.3e-17, 0.705, 0.981 | PDLC01440,Csm5, 2, 2800, 0.023, 0.04 | PDLC01441,COG1336, 1, 11, 0.032, 0.073 | PDLC01441,COG1336, 2, 0.024, 0.036, 0.082 | PDLC01442,COG1337, 1, 2.2e-05, 0.061, 0.115 | PDLC01571,mkCas0182, 1, 3.4e-16, 0.358, 0.552 | PDLC01571,mkCas0182, 2, 13, 0.116, 0.133 | PDLC01613,pfam03787, 1, 1.3e-08, 0.279, 0.288 | PDLC01733,COG1332, 1, 4.5e-11, 0.358, 0.501 | PDLC01733,COG1332, 2, 280, 0.143, 0.225 | PDLC01733,COG1332, 3, 480, 0.045, 0.068","PDLC01440, Csm5, 1.3e-17, 0.705, 0.981 | PDLC01571, mkCas0182, 3.4e-16, 0.358, 0.552 | PDLC01275, cd09662, 2.5e-12, 0.358, 0.52 | PDLC01733, COG1332, 4.5e-11, 0.358, 0.501 | PDLC01020, cas_TM1807_csm5, 6.5e-10, 0.175, 0.258"
3,NZ_CP025084.1,cas_type_III-A,WP_021014789.1,PDLC02098,Cas6_IIIa_Cas6_IIIa,Cas6_IIIa,4.5999999999999994e-42,5.1999999999999994e-42,0.958,0.99,4383055,4383978,+,CRISPR system precrRNA processing endoribonuclease RAMP protein Cas6 [Serratia sp. ATCC 39006],3850,4398,"PDLC01373,cd09760, 1, 0.00032, 0.248, 0.256 | PDLC01373,cd09760, 2, 140, 0.179, 0.187 | PDLC01373,cd09760, 3, 980, 0.072, 0.076 | PDLC01466,COG5551, 1, 0.00022, 0.443, 0.538 | PDLC01477,mkCas0066, 1, 1.6e-92, 0.967, 0.983 | PDLC01496,mkCas0091, 1, 5.7e-91, 0.984, 0.989 | PDLC01650,pfam10040, 1, 5.9e-19, 0.375, 0.99 | PDLC02098,Cas6_IIIa_Cas6_IIIa, 1, 5.2e-42, 0.958, 0.99","PDLC01477, mkCas0066, 1.6e-92, 0.967, 0.983 | PDLC01496, mkCas0091, 5.7e-91, 0.984, 0.989 | PDLC02098, Cas6_IIIa_Cas6_IIIa, 5.2e-42, 0.958, 0.99 | PDLC01650, pfam10040, 5.9e-19, 0.375, 0.99 | PDLC01466, COG5551, 0.00022, 0.443, 0.538"
3,NZ_CP025084.1,cas_type_III-A,WP_021014788.1,PDLC01051,shah_acc_0045,NucC,6.199999999999998e-96,6.899999999999998e-96,0.984,0.984,4384031,4384783,-,hypothetical protein [Serratia sp. ATCC 39006],3851,4398,"PDLC01051,shah_acc_0045, 1, 6.9e-96, 0.984, 0.984 | PDLC01495,mkCas0090, 1, 1.1e-36, 0.476, 0.967","PDLC01051, shah_acc_0045, 6.9e-96, 0.984, 0.984 | PDLC01495, mkCas0090, 1.1e-36, 0.476, 0.967"
4,NZ_CP025084.1,CRISPR_array,CRISPR004,NA,NA,CRISPR_array,NA,6.2,NA,NA,4385117,4385714,+,CRISPR004; repeat=GTCCGTAAGGACGTTCCCTGACTGAAGGGATTAAGAC; score=6.20,3851.04,4398,NA,NA
1,NZ_CP025084.1,AbiE,WP_021014005.1,PDLC02296,AbiEii_WP_066409903.1,AbiEii,3.6999999999999987e-104,4.0999999999999986e-104,0.946,0.965,243531,244418,-,nucleotidyl transferase AbiEii/AbiGii toxin family protein [Serratia sp. ATCC 39006],215,4398,"PDLC02289,AbiEii_WP_007349585.1, 1, 4.9e-06, 0.251, 0.252 | PDLC02289,AbiEii_WP_007349585.1, 2, 24, 0.197, 0.194 | PDLC02291,AbiEii_WP_082807810.1, 1, 5.8e-07, 0.546, 0.49 | PDLC02291,AbiEii_WP_082807810.1, 2, 100, 0.156, 0.142 | PDLC02292,AbiEii_WP_010527912.1, 1, 4.8e-05, 0.251, 0.244 | PDLC02292,AbiEii_WP_010527912.1, 2, 0.012, 0.325, 0.357 | PDLC02293,AbiEii_WP_045959881.1, 1, 1.5e-17, 0.827, 0.885 | PDLC02294,AbiEii_WP_099148274.1, 1, 1.3e-06, 0.783, 0.827 | PDLC02296,AbiEii_WP_066409903.1, 1, 4.1e-104, 0.946, 0.965 | PDLC02297,AbiEii_WP_106546964.1, 1, 9.6e-05, 0.559, 0.573 | PDLC02298,AbiEii_WP_085578968.1, 1, 0.29, 0.085, 0.114 | PDLC02298,AbiEii_WP_085578968.1, 2, 0.00072, 0.322, 0.409 | PDLC02299,AbiEii_WP_105958957.1, 1, 0.0068, 0.553, 0.448 | PDLC02302,AbiEii_WP_076406552.1, 1, 9.6e-08, 0.563, 0.562 | PDLC02303,AbiEii_WP_111872158.1, 1, 1.5e-06, 0.559, 0.61 | PDLC02304,AbiEii_WP_034042188.1, 1, 2.9e-22, 0.739, 0.812 | PDLC02305,AbiEii_WP_096461967.1, 1, 1e-05, 0.614, 0.569 | PDLC02306,AbiEii_WP_084590683.1, 1, 1.3e-06, 0.559, 0.625 | PDLC02306,AbiEii_WP_084590683.1, 2, 120, 0.132, 0.139 | PDLC02307,AbiEii_WP_156423273.1, 1, 2.1e-11, 0.766, 0.881 | PDLC02313,AbiEii_WP_099005948.1, 1, 4.1e-15, 0.298, 0.35 | PDLC02313,AbiEii_WP_099005948.1, 2, 0.079, 0.247, 0.264 | PDLC02317,AbiEii_WP_096360271.1, 1, 3.9e-10, 0.644, 0.495 | PDLC02318,AbiEii_WP_069691453.1, 1, 2.3e-12, 0.607, 0.596 | PDLC02321,AbiEii_WP_169730291.1, 1, 0.0029, 0.159, 0.159 | PDLC02321,AbiEii_WP_169730291.1, 2, 0.00028, 0.244, 0.243 | PDLC02323,AbiEii_WP_077075795.1, 1, 1.3e-17, 0.79, 0.863 | PDLC02324,AbiEii_WP_084488417.1, 1, 0.00049, 0.122, 0.156 | PDLC02324,AbiEii_WP_084488417.1, 2, 2.8e-06, 0.308, 0.372 | PDLC02328,AbiEii_WP_009233131.1, 1, 9.5e-07, 0.719, 0.882 | PDLC02330,AbiEii_WP_028841950.1, 1, 1.1e-14, 0.79, 0.954","PDLC02296, AbiEii_WP_066409903.1, 4.1e-104, 0.946, 0.965 | PDLC02304, AbiEii_WP_034042188.1, 2.9e-22, 0.739, 0.812 | PDLC02323, AbiEii_WP_077075795.1, 1.3e-17, 0.79, 0.863 | PDLC02293, AbiEii_WP_045959881.1, 1.5e-17, 0.827, 0.885 | PDLC02313, AbiEii_WP_099005948.1, 4.1e-15, 0.298, 0.35"
1,NZ_CP025084.1,AbiE,WP_021014004.1,PDLC02232,AbiEi_WP_050009329.1,AbiEi,1.7999999999999998e-62,1.9999999999999996e-62,0.977,0.949,244447,244971,-,DUF4095 domain-containing protein [Serratia sp. ATCC 39006],216,4398,"PDLC02226,AbiEi_WP_146016717.1, 1, 0.038, 0.144, 0.124 | PDLC02230,AbiEi_WP_022933255.1, 1, 9.6e-07, 0.678, 0.573 | PDLC02232,AbiEi_WP_050009329.1, 1, 2e-62, 0.977, 0.949 | PDLC02240,AbiEi_WP_013606017.1, 1, 0.00096, 0.5, 0.398 | PDLC02241,AbiEi_WP_139786902.1, 1, 4e-07, 0.546, 0.452 | PDLC02256,AbiEi_WP_102372703.1, 1, 0.014, 0.42, 0.402 | PDLC02265,AbiEi_WP_076488363.1, 1, 0.0061, 0.276, 0.242 | PDLC02267,AbiEi_WP_082871982.1, 1, 0.00052, 0.649, 0.425 | PDLC02272,AbiEi_WP_005862062.1, 1, 1.1e-06, 0.534, 0.445 | PDLC02274,AbiEi_WP_020504080.1, 1, 0.00036, 0.46, 0.359 | PDLC02275,AbiEi_WP_006905458.1, 1, 0.0041, 0.316, 0.293 | PDLC02283,AbiEi_pseudo_subWP_007706639.1, 1, 0.0053, 0.282, 0.244 | PDLC02283,AbiEi_pseudo_subWP_007706639.1, 2, 520, 0.098, 0.085","PDLC02232, AbiEi_WP_050009329.1, 2e-62, 0.977, 0.949 | PDLC02241, AbiEi_WP_139786902.1, 4e-07, 0.546, 0.452 | PDLC02230, AbiEi_WP_022933255.1, 9.6e-07, 0.678, 0.573 | PDLC02272, AbiEi_WP_005862062.1, 1.1e-06, 0.534, 0.445 | PDLC02274, AbiEi_WP_020504080.1, 0.00036, 0.46, 0.359"
2,NZ_CP025084.1,AbiE,WP_021013440.1,PDLC02290,AbiEii_WP_067065479.1,AbiEii,8.499999999999999e-121,9.799999999999997e-121,0.967,0.986,923883,924800,-,nucleotidyl transferase AbiEii/AbiGii toxin family protein [Serratia sp. ATCC 39006],811,4398,"PDLC02288,AbiEii_WP_110023304.1, 1, 0.0032, 0.239, 0.231 | PDLC02288,AbiEii_WP_110023304.1, 2, 0.39, 0.069, 0.071 | PDLC02289,AbiEii_WP_007349585.1, 1, 0.069, 0.393, 0.411 | PDLC02290,AbiEii_WP_067065479.1, 1, 9.8e-121, 0.967, 0.986 | PDLC02291,AbiEii_WP_082807810.1, 1, 1.2e-06, 0.515, 0.503 | PDLC02291,AbiEii_WP_082807810.1, 2, 190, 0.095, 0.09 | PDLC02292,AbiEii_WP_010527912.1, 1, 0.014, 0.367, 0.371 | PDLC02292,AbiEii_WP_010527912.1, 2, 0.66, 0.115, 0.102 | PDLC02293,AbiEii_WP_045959881.1, 1, 0.00028, 0.469, 0.548 | PDLC02294,AbiEii_WP_099148274.1, 1, 2.6e-12, 0.528, 0.612 | PDLC02295,AbiEii_HBX79544.1, 1, 0.083, 0.138, 0.146 | PDLC02298,AbiEii_WP_085578968.1, 1, 8.8e-07, 0.489, 0.623 | PDLC02299,AbiEii_WP_105958957.1, 1, 0.00022, 0.105, 0.093 | PDLC02303,AbiEii_WP_111872158.1, 1, 5.8e-13, 0.515, 0.618 | PDLC02304,AbiEii_WP_034042188.1, 1, 2e-13, 0.544, 0.642 | PDLC02304,AbiEii_WP_034042188.1, 2, 1400, 0.026, 0.031 | PDLC02305,AbiEii_WP_096461967.1, 1, 6e-31, 0.833, 0.853 | PDLC02307,AbiEii_WP_156423273.1, 1, 1e-07, 0.528, 0.626 | PDLC02313,AbiEii_WP_099005948.1, 1, 8.8e-05, 0.479, 0.579 | PDLC02316,AbiEii_WP_074501794.1, 1, 0.098, 0.134, 0.131 | PDLC02316,AbiEii_WP_074501794.1, 2, 400, 0.118, 0.137 | PDLC02317,AbiEii_WP_096360271.1, 1, 50, 0.187, 0.139 | PDLC02317,AbiEii_WP_096360271.1, 2, 0.019, 0.216, 0.167 | PDLC02318,AbiEii_WP_069691453.1, 1, 45, 0.069, 0.075 | PDLC02318,AbiEii_WP_069691453.1, 2, 4.2e-07, 0.508, 0.539 | PDLC02323,AbiEii_WP_077075795.1, 1, 0.00027, 0.528, 0.645 | PDLC02324,AbiEii_WP_084488417.1, 1, 4.8e-09, 0.485, 0.571 | PDLC02326,AbiEii_WP_096298108.1, 1, 0.25, 0.131, 0.301 | PDLC02326,AbiEii_WP_096298108.1, 2, 110, 0.108, 0.248 | PDLC02328,AbiEii_WP_009233131.1, 1, 1.7e-06, 0.489, 0.65 | PDLC02330,AbiEii_WP_028841950.1, 1, 0.0071, 0.485, 0.616","PDLC02290, AbiEii_WP_067065479.1, 9.8e-121, 0.967, 0.986 | PDLC02305, AbiEii_WP_096461967.1, 6e-31, 0.833, 0.853 | PDLC02304, AbiEii_WP_034042188.1, 2e-13, 0.544, 0.642 | PDLC02303, AbiEii_WP_111872158.1, 5.8e-13, 0.515, 0.618 | PDLC02294, AbiEii_WP_099148274.1, 2.6e-12, 0.528, 0.612"
2,NZ_CP025084.1,AbiE,WP_037380309.1,PDLC02227,AbiEi_WP_068866247.1,AbiEi,2.4999999999999993e-82,2.799999999999999e-82,0.965,0.97,924793,925566,-,type IV toxin-antitoxin system AbiEi family antitoxin [Serratia sp. ATCC 39006],812,4398,"PDLC02225,AbiEi_WP_047105540.1, 1, 0.019, 0.21, 0.263 | PDLC02227,AbiEi_WP_068866247.1, 1, 2.8e-82, 0.965, 0.97","PDLC02227, AbiEi_WP_068866247.1, 2.8e-82, 0.965, 0.97 | PDLC02225, AbiEi_WP_047105540.1, 0.019, 0.21, 0.263"
3,NZ_CP025084.1,AbiE,WP_021017652.1,PDLC02232,AbiEi_WP_050009329.1,AbiEi,8.499999999999999e-78,9.5e-78,0.989,0.989,1451617,1452156,+,DUF6088 family protein [Serratia sp. ATCC 39006],1274,4398,"PDLC02225,AbiEi_WP_047105540.1, 1, 7.3e-08, 0.52, 0.414 | PDLC02226,AbiEi_WP_146016717.1, 1, 1.8e-10, 0.642, 0.554 | PDLC02227,AbiEi_WP_068866247.1, 1, 0.022, 0.447, 0.318 | PDLC02228,AbiEi_OGS01369.1, 1, 1.7e-05, 0.385, 0.301 | PDLC02229,AbiEi_WP_092960020.1, 1, 0.006, 0.324, 0.42 | PDLC02230,AbiEi_WP_022933255.1, 1, 2.1e-11, 0.687, 0.599 | PDLC02232,AbiEi_WP_050009329.1, 1, 9.5e-78, 0.989, 0.989 | PDLC02233,AbiEi_WP_060913257.1, 1, 0.0066, 0.631, 0.533 | PDLC02235,AbiEi_WP_103474522.1, 1, 0.0043, 0.235, 0.192 | PDLC02236,AbiEi_WP_025580240.1, 1, 0.0059, 0.419, 0.391 | PDLC02240,AbiEi_WP_013606017.1, 1, 6.7e-08, 0.626, 0.505 | PDLC02241,AbiEi_WP_139786902.1, 1, 2.3e-13, 0.754, 0.623 | PDLC02247,AbiEi_WP_023355414.1, 1, 3.1e-05, 0.486, 0.405 | PDLC02248,AbiEi_WP_014757546.1, 1, 200, 0.207, 0.172 | PDLC02248,AbiEi_WP_014757546.1, 2, 0.016, 0.553, 0.47 | PDLC02249,AbiEi_NJD28597.1, 1, 0.00011, 0.726, 0.641 | PDLC02255,AbiEi_WP_026161743.1, 1, 3.9e-06, 0.542, 0.468 | PDLC02260,AbiEi_WP_157044108.1, 1, 0.0053, 0.587, 0.74 | PDLC02264,AbiEi_WP_007349584.1, 1, 8.1e-05, 0.62, 0.551 | PDLC02265,AbiEi_WP_076488363.1, 1, 2.5e-06, 0.43, 0.369 | PDLC02266,AbiEi_WP_170110179.1, 1, 1.8e-10, 0.754, 0.527 | PDLC02267,AbiEi_WP_082871982.1, 1, 5e-14, 0.715, 0.468 | PDLC02269,AbiEi_WP_101304315.1, 1, 0.00036, 0.48, 0.327 | PDLC02270,AbiEi_WP_019177799.1, 1, 0.0037, 0.637, 0.43 | PDLC02272,AbiEi_WP_005862062.1, 1, 9.7e-09, 0.631, 0.52 | PDLC02274,AbiEi_WP_020504080.1, 1, 4.6e-08, 0.587, 0.461 | PDLC02275,AbiEi_WP_006905458.1, 1, 0.013, 0.48, 0.44 | PDLC02276,AbiEi_WP_069691454.1, 1, 0.00022, 0.587, 0.381 | PDLC02282,AbiEi_WP_069175104.1, 1, 1.4e-08, 0.726, 0.504 | PDLC02283,AbiEi_pseudo_subWP_007706639.1, 1, 2.4e-05, 0.397, 0.333 | PDLC02287,AbiEi_WP_009249990.1, 1, 0.0011, 0.631, 0.419","PDLC02232, AbiEi_WP_050009329.1, 9.5e-78, 0.989, 0.989 | PDLC02267, AbiEi_WP_082871982.1, 5e-14, 0.715, 0.468 | PDLC02241, AbiEi_WP_139786902.1, 2.3e-13, 0.754, 0.623 | PDLC02230, AbiEi_WP_022933255.1, 2.1e-11, 0.687, 0.599 | PDLC02226, AbiEi_WP_146016717.1, 1.8e-10, 0.642, 0.554 | PDLC02266, AbiEi_WP_170110179.1, 1.8e-10, 0.754, 0.527"
3,NZ_CP025084.1,AbiE,WP_021017651.1,PDLC02296,AbiEii_WP_066409903.1,AbiEii,5.499999999999999e-123,6.3e-123,0.938,0.986,1452146,1453069,+,nucleotidyl transferase AbiEii/AbiGii toxin family protein [Serratia sp. ATCC 39006],1275,4398,"PDLC02289,AbiEii_WP_007349585.1, 1, 1.1e-07, 0.306, 0.282 | PDLC02289,AbiEii_WP_007349585.1, 2, 370, 0.072, 0.058 | PDLC02291,AbiEii_WP_082807810.1, 1, 3.4e-09, 0.55, 0.487 | PDLC02292,AbiEii_WP_010527912.1, 1, 3.6e-11, 0.375, 0.36 | PDLC02293,AbiEii_WP_045959881.1, 1, 2.2e-22, 0.765, 0.841 | PDLC02294,AbiEii_WP_099148274.1, 1, 8e-08, 0.779, 0.85 | PDLC02295,AbiEii_HBX79544.1, 1, 0.0043, 0.564, 0.632 | PDLC02296,AbiEii_WP_066409903.1, 1, 6.3e-123, 0.938, 0.986 | PDLC02297,AbiEii_WP_106546964.1, 1, 3.6e-07, 0.541, 0.554 | PDLC02298,AbiEii_WP_085578968.1, 1, 0.0064, 0.642, 0.75 | PDLC02299,AbiEii_WP_105958957.1, 1, 0.0017, 0.537, 0.433 | PDLC02302,AbiEii_WP_076406552.1, 1, 2.6e-08, 0.596, 0.594 | PDLC02303,AbiEii_WP_111872158.1, 1, 0.0081, 0.534, 0.578 | PDLC02304,AbiEii_WP_034042188.1, 1, 2.1e-20, 0.648, 0.7 | PDLC02306,AbiEii_WP_084590683.1, 1, 3.2e-05, 0.56, 0.625 | PDLC02307,AbiEii_WP_156423273.1, 1, 1.1e-07, 0.101, 0.119 | PDLC02307,AbiEii_WP_156423273.1, 2, 1.5, 0.228, 0.301 | PDLC02313,AbiEii_WP_099005948.1, 1, 8.5e-15, 0.733, 0.807 | PDLC02315,AbiEii_WP_110076847.1, 1, 0.00011, 0.218, 0.199 | PDLC02316,AbiEii_WP_074501794.1, 1, 0.0045, 0.238, 0.229 | PDLC02317,AbiEii_WP_096360271.1, 1, 1e-08, 0.616, 0.475 | PDLC02318,AbiEii_WP_069691453.1, 1, 2.8e-14, 0.609, 0.593 | PDLC02319,AbiEii_WP_148235064.1, 1, 4.7e-05, 0.56, 0.647 | PDLC02321,AbiEii_WP_169730291.1, 1, 2.6e-05, 0.156, 0.162 | PDLC02321,AbiEii_WP_169730291.1, 2, 0.0024, 0.414, 0.402 | PDLC02322,AbiEii_WP_066910913.1, 1, 8.1e-06, 0.254, 0.231 | PDLC02323,AbiEii_WP_077075795.1, 1, 5.1e-18, 0.759, 0.847 | PDLC02324,AbiEii_WP_084488417.1, 1, 0.00044, 0.101, 0.134 | PDLC02324,AbiEii_WP_084488417.1, 2, 0.0076, 0.3, 0.407 | PDLC02327,AbiEii_WP_052604370.1, 1, 0.021, 0.107, 0.205 | PDLC02328,AbiEii_WP_009233131.1, 1, 1.2e-08, 0.616, 0.754 | PDLC02330,AbiEii_WP_028841950.1, 1, 9.1e-13, 0.179, 0.251 | PDLC02330,AbiEii_WP_028841950.1, 2, 0.21, 0.192, 0.256","PDLC02296, AbiEii_WP_066409903.1, 6.3e-123, 0.938, 0.986 | PDLC02293, AbiEii_WP_045959881.1, 2.2e-22, 0.765, 0.841 | PDLC02304, AbiEii_WP_034042188.1, 2.1e-20, 0.648, 0.7 | PDLC02323, AbiEii_WP_077075795.1, 5.1e-18, 0.759, 0.847 | PDLC02313, AbiEii_WP_099005948.1, 8.5e-15, 0.733, 0.807"
2,NZ_CP025084.1,RM_type_I,WP_021014229.1,PDLC03019,MTase_I_00002,MTase_I,5.199999999999999e-174,5.799999999999999e-172,0.979,0.534,21859,23565,+,type I restriction-modification system subunit M [Serratia sp. ATCC 39006],21,4398,"PDLC03018,MTase_I_00001, 1, 3.3e-09, 0.13, 0.096 | PDLC03018,MTase_I_00001, 2, 0.021, 0.1, 0.076 | PDLC03019,MTase_I_00002, 1, 5.8e-172, 0.979, 0.534 | PDLC03020,MTase_I_00003, 1, 2.9e-06, 0.079, 0.11 | PDLC03020,MTase_I_00003, 2, 2.2e-31, 0.393, 0.563 | PDLC03021,MTase_I_00004, 1, 7.1e-52, 0.824, 0.894 | PDLC03022,MTase_I_00005, 1, 2.9e-83, 0.914, 0.559 | PDLC03025,MTase_I_00008, 1, 8.5e-24, 0.496, 0.473 | PDLC03026,MTase_I_00009, 1, 19, 0.067, 0.08 | PDLC03026,MTase_I_00009, 2, 3.8e-37, 0.569, 0.655 | PDLC03027,MTase_I_00010, 1, 1.9e-10, 0.088, 0.062 | PDLC03027,MTase_I_00010, 2, 1.2e-57, 0.627, 0.411 | PDLC03028,MTase_I_00011, 1, 5.1e-05, 0.088, 0.04 | PDLC03028,MTase_I_00011, 2, 3.9e-48, 0.641, 0.293 | PDLC03029,MTase_I_00012, 1, 0.0029, 0.095, 0.082 | PDLC03029,MTase_I_00012, 2, 8.6e-48, 0.563, 0.492 | PDLC03030,MTase_I_00013, 1, 2.4e-05, 0.257, 0.237 | PDLC03031,MTase_I_00014, 1, 1.9e-81, 0.924, 0.591 | PDLC03032,MTase_I_00015, 1, 7.8e-08, 0.07, 0.04 | PDLC03032,MTase_I_00015, 2, 8.5e-35, 0.592, 0.318 | PDLC03033,MTase_I_00016, 1, 4.7e-32, 0.699, 0.715 | PDLC03034,MTase_I_00017, 1, 2.8e-06, 0.116, 0.095 | PDLC03034,MTase_I_00017, 2, 2.6, 0.174, 0.149 | PDLC03035,MTase_I_00018, 1, 7.5e-85, 0.833, 0.643 | PDLC03035,MTase_I_00018, 2, 1.5e-15, 0.136, 0.118 | PDLC03036,MTase_I_00019, 1, 1.8e-15, 0.394, 0.354 | PDLC03037,MTase_I_00020, 1, 1.5e-28, 0.424, 0.292 | PDLC03037,MTase_I_00020, 2, 0.57, 0.1, 0.076 | PDLC03038,MTase_I_00021, 1, 0.00026, 0.083, 0.052 | PDLC03038,MTase_I_00021, 2, 7.8e-50, 0.692, 0.417 | PDLC03039,MTase_I_00022, 1, 3e-42, 0.905, 0.633","PDLC03019, MTase_I_00002, 5.8e-172, 0.979, 0.534 | PDLC03035, MTase_I_00018, 7.5e-85, 0.833, 0.643 | PDLC03022, MTase_I_00005, 2.9e-83, 0.914, 0.559 | PDLC03031, MTase_I_00014, 1.9e-81, 0.924, 0.591 | PDLC03027, MTase_I_00010, 1.2e-57, 0.627, 0.411"
2,NZ_CP025084.1,RM_type_I,WP_021014228.1,PDLC03099,Specificity_I_00048,Specificity_I,4.9999999999999987e-138,5.599999999999999e-138,0.998,0.998,23555,24877,+,restriction endonuclease subunit S [Serratia sp. ATCC 39006],22,4398,"PDLC03019,MTase_I_00002, 1, 1.4e-06, 0.168, 0.078 | PDLC03019,MTase_I_00002, 2, 0.096, 0.089, 0.041 | PDLC03019,MTase_I_00002, 3, 6.6e-08, 0.123, 0.058 | PDLC03032,MTase_I_00015, 1, 140, 0.223, 0.103 | PDLC03032,MTase_I_00015, 2, 0.0035, 0.198, 0.085 | PDLC03038,MTase_I_00021, 1, 0.0078, 0.275, 0.137 | PDLC03052,Specificity_I_00001, 1, 1.1e-29, 0.323, 0.306 | PDLC03052,Specificity_I_00001, 2, 4.6e-06, 0.195, 0.185 | PDLC03054,Specificity_I_00003, 1, 4.1e-32, 0.364, 0.394 | PDLC03054,Specificity_I_00003, 2, 0.81, 0.048, 0.052 | PDLC03055,Specificity_I_00004, 1, 0.0028, 0.168, 0.192 | PDLC03055,Specificity_I_00004, 2, 0.22, 0.075, 0.082 | PDLC03058,Specificity_I_00007, 1, 210, 0.082, 0.092 | PDLC03058,Specificity_I_00007, 2, 0.0046, 0.293, 0.341 | PDLC03059,Specificity_I_00008, 1, 7.5e-05, 0.364, 0.408 | PDLC03059,Specificity_I_00008, 2, 120, 0.059, 0.063 | PDLC03061,Specificity_I_00010, 1, 3.1e-20, 0.316, 0.389 | PDLC03061,Specificity_I_00010, 2, 23, 0.164, 0.197 | PDLC03062,Specificity_I_00011, 1, 0.0032, 0.195, 0.208 | PDLC03062,Specificity_I_00011, 2, 0.52, 0.402, 0.485 | PDLC03063,Specificity_I_00012, 1, 1.3e-63, 0.402, 0.474 | PDLC03063,Specificity_I_00012, 2, 1.6e-11, 0.477, 0.575 | PDLC03064,Specificity_I_00013, 1, 6.3e-05, 0.318, 0.342 | PDLC03064,Specificity_I_00013, 2, 36, 0.191, 0.203 | PDLC03065,Specificity_I_00014, 1, 7.2e-18, 0.282, 0.347 | PDLC03065,Specificity_I_00014, 2, 180, 0.084, 0.102 | PDLC03065,Specificity_I_00014, 3, 2.6e-08, 0.189, 0.231 | PDLC03066,Specificity_I_00015, 1, 2.1e-41, 0.773, 0.701 | PDLC03068,Specificity_I_00017, 1, 6.4e-24, 0.282, 0.315 | PDLC03068,Specificity_I_00017, 2, 1.3e-57, 0.775, 0.725 | PDLC03069,Specificity_I_00018, 1, 4.6, 0.15, 0.168 | PDLC03069,Specificity_I_00018, 2, 7.7e-09, 0.284, 0.336 | PDLC03072,Specificity_I_00021, 1, 1.2e-05, 0.207, 0.223 | PDLC03072,Specificity_I_00021, 2, 0.0038, 0.443, 0.478 | PDLC03073,Specificity_I_00022, 1, 1.4e-05, 0.216, 0.233 | PDLC03073,Specificity_I_00022, 2, 1, 0.191, 0.19 | PDLC03074,Specificity_I_00023, 1, 1.1e-09, 0.255, 0.277 | PDLC03074,Specificity_I_00023, 2, 2.5e-14, 0.432, 0.475 | PDLC03075,Specificity_I_00024, 1, 0.041, 0.159, 0.174 | PDLC03075,Specificity_I_00024, 2, 4.9, 0.057, 0.061 | PDLC03078,Specificity_I_00027, 1, 7.1e-05, 0.336, 0.415 | PDLC03078,Specificity_I_00027, 2, 200, 0.07, 0.076 | PDLC03079,Specificity_I_00028, 1, 2.1e-09, 0.864, 0.779 | PDLC03082,Specificity_I_00031, 1, 3.9e-36, 0.77, 0.905 | PDLC03083,Specificity_I_00032, 1, 1.9e-12, 0.436, 0.271 | PDLC03084,Specificity_I_00033, 1, 640, 0.045, 0.051 | PDLC03084,Specificity_I_00033, 2, 0.00046, 0.2, 0.232 | PDLC03084,Specificity_I_00033, 3, 8.9, 0.218, 0.253 | PDLC03086,Specificity_I_00035, 1, 75, 0.052, 0.05 | PDLC03086,Specificity_I_00035, 2, 1e-81, 0.877, 0.834 | PDLC03087,Specificity_I_00036, 1, 2.6e-07, 0.257, 0.289 | PDLC03087,Specificity_I_00036, 2, 8e-06, 0.432, 0.486 | PDLC03088,Specificity_I_00037, 1, 350, 0.184, 0.134 | PDLC03088,Specificity_I_00037, 2, 3.5e-07, 0.35, 0.239 | PDLC03089,Specificity_I_00038, 1, 4.2e-101, 0.991, 0.996 | PDLC03090,Specificity_I_00039, 1, 9.4e-07, 0.245, 0.253 | PDLC03090,Specificity_I_00039, 2, 6.8e-05, 0.314, 0.339 | PDLC03090,Specificity_I_00039, 3, 33, 0.061, 0.062 | PDLC03092,Specificity_I_00041, 1, 3.7e-61, 0.95, 0.977 | PDLC03093,Specificity_I_00042, 1, 5.8e-09, 0.309, 0.358 | PDLC03096,Specificity_I_00045, 1, 1.6, 0.152, 0.111 | PDLC03096,Specificity_I_00045, 2, 0.00093, 0.22, 0.153 | PDLC03098,Specificity_I_00047, 1, 5.8e-10, 0.361, 0.4 | PDLC03098,Specificity_I_00047, 2, 3.3e-07, 0.445, 0.454 | PDLC03099,Specificity_I_00048, 1, 5.6e-138, 0.998, 0.998 | PDLC03100,Specificity_I_00049, 1, 2.8e-05, 0.275, 0.332 | PDLC03100,Specificity_I_00049, 2, 2.6e-11, 0.293, 0.332 | PDLC03101,Specificity_I_00050, 1, 4.3e-07, 0.314, 0.397 | PDLC03101,Specificity_I_00050, 2, 0.1, 0.289, 0.338 | PDLC03102,Specificity_I_00051, 1, 6.8e-22, 0.375, 0.428 | PDLC03103,Specificity_I_00052, 1, 3.1, 0.205, 0.24 | PDLC03103,Specificity_I_00052, 2, 0.018, 0.348, 0.395 | PDLC03104,Specificity_I_00053, 1, 2.9e-11, 0.32, 0.354 | PDLC03104,Specificity_I_00053, 2, 17, 0.118, 0.123 | PDLC03104,Specificity_I_00053, 3, 0.0019, 0.175, 0.186 | PDLC03105,Specificity_I_00054, 1, 0.0034, 0.236, 0.246 | PDLC03105,Specificity_I_00054, 2, 9.5e-09, 0.414, 0.442 | PDLC03106,Specificity_I_00055, 1, 0.12, 0.166, 0.156 | PDLC03106,Specificity_I_00055, 2, 23, 0.048, 0.048 | PDLC03108,Specificity_I_00057, 1, 3.6e-13, 0.775, 0.662 | PDLC03112,Specificity_I_00061, 1, 8.5e-13, 0.193, 0.23 | PDLC03112,Specificity_I_00061, 2, 170, 0.093, 0.106 | PDLC03112,Specificity_I_00061, 3, 150, 0.073, 0.085 | PDLC03112,Specificity_I_00061, 4, 0.0011, 0.107, 0.124 | PDLC03113,Specificity_I_00062, 1, 0.0045, 0.209, 0.225 | PDLC03113,Specificity_I_00062, 2, 0.11, 0.416, 0.469 | PDLC03115,Specificity_I_00064, 1, 6.3e-18, 0.314, 0.294 | PDLC03116,Specificity_I_00065, 1, 1.4e-36, 0.314, 0.335 | PDLC03116,Specificity_I_00065, 2, 16, 0.045, 0.049 | PDLC03119,Specificity_I_00068, 1, 8.2e-06, 0.227, 0.26 | PDLC03119,Specificity_I_00068, 2, 62, 0.059, 0.064 | PDLC03119,Specificity_I_00068, 3, 25, 0.175, 0.193 | PDLC03121,Specificity_I_00070, 1, 0.082, 0.107, 0.116 | PDLC03121,Specificity_I_00070, 2, 0.0068, 0.2, 0.224 | PDLC03123,Specificity_I_00072, 1, 0.0093, 0.184, 0.195 | PDLC03123,Specificity_I_00072, 2, 0.012, 0.066, 0.072 | PDLC03124,Specificity_I_00073, 1, 2.8e-06, 0.377, 0.448 | PDLC03124,Specificity_I_00073, 2, 10, 0.218, 0.235 | PDLC03126,Specificity_I_00075, 1, 1, 0.125, 0.084 | PDLC03126,Specificity_I_00075, 2, 1.1e-19, 0.266, 0.177 | PDLC03127,Specificity_I_00076, 1, 71, 0.052, 0.476 | PDLC03127,Specificity_I_00076, 2, 0.00032, 0.289, 0.242 | PDLC03130,Specificity_I_00079, 1, 1.3e-23, 0.33, 0.308 | PDLC03130,Specificity_I_00079, 2, 3.6e-31, 0.286, 0.29 | PDLC03130,Specificity_I_00079, 3, 0.015, 0.102, 0.102 | PDLC03132,Specificity_I_00081, 1, 1.3e-06, 0.186, 0.196 | PDLC03132,Specificity_I_00081, 2, 930, 0.034, 0.039 | PDLC03132,Specificity_I_00081, 3, 0.00051, 0.134, 0.152 | PDLC03133,Specificity_I_00082, 1, 7.6e-05, 0.159, 0.165 | PDLC03133,Specificity_I_00082, 2, 0.021, 0.166, 0.175 | PDLC03134,Specificity_I_00083, 1, 250, 0.07, 0.077 | PDLC03134,Specificity_I_00083, 2, 6.5e-06, 0.173, 0.182 | PDLC03134,Specificity_I_00083, 3, 7.9, 0.057, 0.058 | PDLC03134,Specificity_I_00083, 4, 0.94, 0.068, 0.07 | PDLC03135,Specificity_I_00084, 1, 1.9e-11, 0.202, 0.155 | PDLC03135,Specificity_I_00084, 2, 5.9e-33, 0.286, 0.213 | PDLC03135,Specificity_I_00084, 3, 0.037, 0.084, 0.062 | PDLC03136,Specificity_I_00085, 1, 3.3e-31, 0.268, 0.37 | PDLC03136,Specificity_I_00085, 2, 1.7e-14, 0.18, 0.241 | PDLC03136,Specificity_I_00085, 3, 6.9e-11, 0.482, 0.623 | PDLC03137,Specificity_I_00086, 1, 4e-15, 0.375, 0.464 | PDLC03137,Specificity_I_00086, 2, 33, 0.061, 0.074 | PDLC03138,Specificity_I_00087, 1, 1.2e-18, 0.425, 0.392 | PDLC03138,Specificity_I_00087, 2, 1.4e-05, 0.448, 0.4 | PDLC03140,Specificity_I_00089, 1, 0.0022, 0.332, 0.356 | PDLC03144,Specificity_I_00093, 1, 3.8e-09, 0.3, 0.356 | PDLC03144,Specificity_I_00093, 2, 0.036, 0.302, 0.325 | PDLC03148,Specificity_I_00097, 1, 1.1, 0.111, 0.108 | PDLC03148,Specificity_I_00097, 2, 0.69, 0.139, 0.135 | PDLC03148,Specificity_I_00097, 3, 3.4, 0.293, 0.296 | PDLC03149,Specificity_I_00098, 1, 0.01, 0.17, 0.195 | PDLC03149,Specificity_I_00098, 2, 0.017, 0.075, 0.082 | PDLC03152,Specificity_I_00101, 1, 0.092, 0.184, 0.206 | PDLC03152,Specificity_I_00101, 2, 4.4e-06, 0.214, 0.233 | PDLC03153,Specificity_I_00102, 1, 0.018, 0.225, 0.249 | PDLC03154,Specificity_I_00103, 1, 1.9e-20, 0.28, 0.313 | PDLC03154,Specificity_I_00103, 2, 8.1e-18, 0.448, 0.522 | PDLC03160,Specificity_I_00109, 1, 1.8e-07, 0.252, 0.28 | PDLC03161,Specificity_I_00110, 1, 9e-07, 0.193, 0.222 | PDLC03161,Specificity_I_00110, 2, 2.3e-07, 0.116, 0.126 | PDLC03162,Specificity_I_00111, 1, 31, 0.1, 0.109 | PDLC03162,Specificity_I_00111, 2, 0.048, 0.223, 0.23 | PDLC03162,Specificity_I_00111, 3, 0.74, 0.064, 0.065 | PDLC03162,Specificity_I_00111, 4, 320, 0.105, 0.107 | PDLC03162,Specificity_I_00111, 5, 170, 0.059, 0.067 | PDLC03163,Specificity_I_00112, 1, 1.4e-08, 0.252, 0.276 | PDLC03163,Specificity_I_00112, 2, 6.3e-07, 0.445, 0.482 | PDLC03164,Specificity_I_00113, 1, 1.7e-09, 0.28, 0.306 | PDLC03164,Specificity_I_00113, 2, 5.6e-12, 0.1, 0.108 | PDLC03164,Specificity_I_00113, 3, 4.7e-22, 0.448, 0.455 | PDLC03165,Specificity_I_00114, 1, 1.8e-08, 0.32, 0.35 | PDLC03165,Specificity_I_00114, 2, 46, 0.177, 0.197 | PDLC03168,Specificity_I_00117, 1, 6.7e-80, 0.993, 0.993 | PDLC03172,Specificity_I_00121, 1, 440, 0.039, 0.039 | PDLC03172,Specificity_I_00121, 2, 1e-07, 0.209, 0.22 | PDLC03172,Specificity_I_00121, 3, 9.9e-20, 0.459, 0.508 | PDLC03177,Specificity_I_00126, 1, 0.15, 0.136, 0.147 | PDLC03177,Specificity_I_00126, 2, 0.00079, 0.077, 0.085 | PDLC03178,Specificity_I_00127, 1, 8.4e-11, 0.361, 0.421 | PDLC03178,Specificity_I_00127, 2, 5.6e-05, 0.43, 0.477 | PDLC03179,Specificity_I_00128, 1, 0.0021, 0.268, 0.216 | PDLC03179,Specificity_I_00128, 2, 5.6e-05, 0.307, 0.248 | PDLC03182,Specificity_I_00131, 1, 0.025, 0.116, 0.114 | PDLC03182,Specificity_I_00131, 2, 400, 0.041, 0.041 | PDLC03182,Specificity_I_00131, 3, 0.12, 0.118, 0.118 | PDLC03184,Specificity_I_00133, 1, 280, 0.182, 0.146 | PDLC03184,Specificity_I_00133, 2, 8.3e-09, 0.425, 0.343 | PDLC03185,Specificity_I_00134, 1, 5.2e-05, 0.241, 0.265 | PDLC03185,Specificity_I_00134, 2, 0.089, 0.341, 0.37 | PDLC03188,Specificity_I_00137, 1, 4.5e-05, 0.245, 0.247 | PDLC03188,Specificity_I_00137, 2, 0.013, 0.259, 0.277 | PDLC03188,Specificity_I_00137, 3, 2.2, 0.055, 0.052 | PDLC03194,Specificity_I_00143, 1, 31, 0.084, 0.102 | PDLC03194,Specificity_I_00143, 2, 12, 0.114, 0.136 | PDLC03194,Specificity_I_00143, 3, 2.2e-13, 0.42, 0.496","PDLC03099, Specificity_I_00048, 5.6e-138, 0.998, 0.998 | PDLC03089, Specificity_I_00038, 4.2e-101, 0.991, 0.996 | PDLC03086, Specificity_I_00035, 1e-81, 0.877, 0.834 | PDLC03168, Specificity_I_00117, 6.7e-80, 0.993, 0.993 | PDLC03063, Specificity_I_00012, 1.3e-63, 0.402, 0.474"
2,NZ_CP025084.1,RM_type_I,WP_021014226.1,PDLC03040,REase_I_00001,REase_I,0,0,0.994,0.989,26058,29192,+,type I restriction endonuclease subunit R [Serratia sp. ATCC 39006],24,4398,"PDLC03040,REase_I_00001, 1, 0, 0.994, 0.989 | PDLC03041,REase_I_00002, 1, 5.6e-10, 0.1, 0.101 | PDLC03041,REase_I_00002, 2, 6.7e-62, 0.473, 0.436 | PDLC03043,REase_I_00004, 1, 2.8e-07, 0.152, 0.505 | PDLC03044,REase_I_00005, 1, 9.3e-51, 0.484, 0.458 | PDLC03044,REase_I_00005, 2, 1.6e-17, 0.08, 0.081 | PDLC03045,REase_I_00006, 1, 0.021, 0.058, 0.063 | PDLC03045,REase_I_00006, 2, 4.5e-10, 0.182, 0.181 | PDLC03045,REase_I_00006, 3, 5.8e-09, 0.081, 0.089 | PDLC03046,REase_I_00007, 1, 6.3e-14, 0.368, 0.38 | PDLC03046,REase_I_00007, 2, 1.5e-13, 0.073, 0.077 | PDLC03048,REase_I_00009, 1, 5.9e-41, 0.424, 0.42 | PDLC03048,REase_I_00009, 2, 7.4e-18, 0.087, 0.092 | PDLC03049,REase_I_00010, 1, 8.6e-07, 0.231, 0.27","PDLC03040, REase_I_00001, 0, 0.994, 0.989 | PDLC03041, REase_I_00002, 6.7e-62, 0.473, 0.436 | PDLC03044, REase_I_00005, 9.3e-51, 0.484, 0.458 | PDLC03048, REase_I_00009, 5.9e-41, 0.424, 0.42 | PDLC03046, REase_I_00007, 6.3e-14, 0.368, 0.38"
1,NZ_CP025084.1,DMS_other,WP_021015404.1,PDLC04135,mads_3,mad3,1.7e-16,1.1e-13,0.943,0.869,3658314,3659795,+,AAA family ATPase [Serratia sp. ATCC 39006],3237,4398,"PDLC02663,DndD_00001, 1, 0.032, 0.043, 0.031 | PDLC02663,DndD_00001, 2, 130, 0.128, 0.093 | PDLC02663,DndD_00001, 3, 0.23, 0.383, 0.271 | PDLC02667,DndD_00005, 1, 0.016, 0.039, 0.029 | PDLC02667,DndD_00005, 2, 5.3, 0.406, 0.289 | PDLC02667,DndD_00005, 3, 2.2, 0.069, 0.05 | PDLC02668,DndD_00006, 1, 0.0025, 0.041, 0.03 | PDLC02668,DndD_00006, 2, 0.0015, 0.556, 0.417 | PDLC02714,PbeC_00006, 1, 0.061, 0.049, 0.037 | PDLC02714,PbeC_00006, 2, 640, 0.041, 0.031 | PDLC02714,PbeC_00006, 3, 5.2, 0.146, 0.114 | PDLC02714,PbeC_00006, 4, 3.6, 0.051, 0.038 | PDLC02740,PbeC_00032, 1, 0.021, 0.041, 0.031 | PDLC02740,PbeC_00032, 2, 0.64, 0.274, 0.208 | PDLC02747,PbeC_00039, 1, 0.0023, 0.065, 0.051 | PDLC02747,PbeC_00039, 2, 61, 0.286, 0.218 | PDLC02756,PbeC_00048, 1, 0.0037, 0.041, 0.031 | PDLC02756,PbeC_00048, 2, 0.065, 0.456, 0.342 | PDLC03660,mREase_IV_00006, 1, 450, 0.032, 0.037 | PDLC03660,mREase_IV_00006, 2, 0.0081, 0.091, 0.104 | PDLC04135,mads_3, 1, 1.1e-13, 0.943, 0.869 | PDLC04140,mads_8, 1, 2.5e-05, 0.86, 0.599","PDLC04135, mads_3, 1.1e-13, 0.943, 0.869 | PDLC04140, mads_8, 2.5e-05, 0.86, 0.599 | PDLC02668, DndD_00006, 0.0015, 0.556, 0.417 | PDLC02747, PbeC_00039, 0.0023, 0.065, 0.051 | PDLC02756, PbeC_00048, 0.0037, 0.041, 0.031"
1,NZ_CP025084.1,DMS_other,pseudo_subWP_076611456.1,PDLC02590,DrmC_00006,DrmC,9.5e-51,1e-50,0.987,0.886,3660940,3661119,+,"transposase, partial [Salmonella enterica]",3240,4398,"PDLC02590,DrmC_00006, 1, 1e-50, 0.987, 0.886 | PDLC04133,mads_1, 1, 440, 0.152, 0.2 | PDLC04133,mads_1, 2, 0.0022, 0.228, 0.3","PDLC02590, DrmC_00006, 1e-50, 0.987, 0.886 | PDLC04133, mads_1, 0.0022, 0.228, 0.3"
3,NZ_CP025084.1,RM_type_IV,WP_021014427.1,PDLC03657,mREase_IV_00003,mREase_IV,1.2999999999999998e-75,1.3999999999999997e-75,0.987,0.984,4775954,4776886,+,restriction endonuclease [Serratia sp. ATCC 39006],4216,4398,"PDLC03657,mREase_IV_00003, 1, 1.4e-75, 0.987, 0.984 | PDLC03663,mREase_IV_00009, 1, 2.4e-10, 0.394, 0.21","PDLC03657, mREase_IV_00003, 1.4e-75, 0.987, 0.984 | PDLC03663, mREase_IV_00009, 2.4e-10, 0.394, 0.21"
2,NZ_CP025084.1,retron_II-A,WP_021017395.1,PDLC02939,retron_II-A1,RT_II-A,9.199999999999998e-110,1.0999999999999997e-109,0.959,0.987,1720550,1721503,-,retron St85 family RNA-directed DNA polymerase [Serratia sp. ATCC 39006],1532,4398,"PDLC02939,retron_II-A1, 1, 1.1e-109, 0.959, 0.987 | PDLC02940,retron_II-A2, 1, 1e-57, 0.89, 0.56 | PDLC02941,retron_II-A3, 1, 5.7e-62, 0.924, 0.896","PDLC02939, retron_II-A1, 1.1e-109, 0.959, 0.987 | PDLC02941, retron_II-A3, 5.7e-62, 0.924, 0.896 | PDLC02940, retron_II-A2, 1e-57, 0.89, 0.56"
2,NZ_CP025084.1,retron_II-A,WP_021017394.1,PDLC02928,retron_type_II_A1_ndt_cluster42_2,NDT_II-A,4e-71,4.699999999999999e-71,0.985,0.982,1721516,1722487,-,retron St85 family effector protein [Serratia sp. ATCC 39006],1533,4398,"PDLC02928,retron_type_II_A1_ndt_cluster42_2, 1, 4.7e-71, 0.985, 0.982 | PDLC02929,retron_type_II_A2_ndt_cluster42_3, 1, 1.4e-06, 0.402, 0.643 | PDLC02929,retron_type_II_A2_ndt_cluster42_3, 2, 480, 0.056, 0.09 | PDLC02930,retron_type_II_A3_ndt_cluster42_1, 1, 2.9e-22, 0.845, 0.853","PDLC02928, retron_type_II_A1_ndt_cluster42_2, 4.7e-71, 0.985, 0.982 | PDLC02930, retron_type_II_A3_ndt_cluster42_1, 2.9e-22, 0.845, 0.853 | PDLC02929, retron_type_II_A2_ndt_cluster42_3, 1.4e-06, 0.402, 0.643"
1,NZ_CP025084.1,retron_I-C,WP_021014561.1,PDLC02966,retron_I-C1,RT-Toprim_I-C,3.199999999999998e-210,3.5999999999999985e-210,0.995,0.965,4625922,4627643,-,retron Ec67 family RNA-directed DNA polymerase/endonuclease [Serratia sp. ATCC 39006],4078,4398,"PDLC02963,retron_type_I_C1_RT_typeIC1, 1, 1.1e-209, 0.993, 0.995 | PDLC02964,retron_type_I_C2_RT_typeIC2, 1, 2.6e-158, 0.983, 0.995 | PDLC02965,retron_type_I_C3_RT_typeIC3, 1, 4e-85, 0.597, 0.626 | PDLC02965,retron_type_I_C3_RT_typeIC3, 2, 0.83, 0.058, 0.059 | PDLC02966,retron_I-C1, 1, 3.6e-210, 0.995, 0.965 | PDLC02967,retron_I-C2, 1, 2.6e-157, 0.981, 0.995 | PDLC02968,retron_I-C3, 1, 2.2e-84, 0.932, 0.957","PDLC02966, retron_I-C1, 3.6e-210, 0.995, 0.965 | PDLC02963, retron_type_I_C1_RT_typeIC1, 1.1e-209, 0.993, 0.995 | PDLC02964, retron_type_I_C2_RT_typeIC2, 2.6e-158, 0.983, 0.995 | PDLC02967, retron_I-C2, 2.6e-157, 0.981, 0.995 | PDLC02965, retron_type_I_C3_RT_typeIC3, 4e-85, 0.597, 0.626"
1,NZ_CP025084.1,retron_I-C,NA,-,TypeIC1_IC2,msr-msd,NA,3.3e-12,NA,NA,4627661,4627793,-,msr-msd identified by match to covariance model: TypeIC1_IC2,4078.011,4398,NA,NA
1,NZ_CP025084.1,Mokosh_TypeII,WP_021014230.1,Mokosh_TypeII__MkoC,Mokosh_TypeII__MkoC,MkoC,1.4999999999999998e-70,2.6999999999999995e-70,0.647,0.615,18263,21550,+,hypothetical protein [Serratia sp. ATCC 39006],20,4398,"Mokosh_TypeII__MkoC,Mokosh_TypeII__MkoC, 1, 2.7e-70, 0.647, 0.615","Mokosh_TypeII__MkoC, Mokosh_TypeII__MkoC, 2.7e-70, 0.647, 0.615"
5,NZ_CP025084.1,SoFic,WP_021014008.1,SoFic__SoFic,SoFic__SoFic,SoFic,2.5999999999999995e-125,2.9999999999999994e-125,0.943,0.97,240323,241426,+,Fic family protein [Serratia sp. ATCC 39006],212,4398,"SoFic__SoFic,SoFic__SoFic, 1, 3e-125, 0.943, 0.97","SoFic__SoFic, SoFic__SoFic, 3e-125, 0.943, 0.97"
4,NZ_CP025084.1,PD-T7-1or5,WP_021016695.1,PD-T7-5_WP_098786838.1,PD-T7-5_WP_098786838.1,PD-T7-5,1.1999999999999998e-116,1.3999999999999997e-116,0.977,0.983,2186733,2187779,-,hypothetical protein [Serratia sp. ATCC 39006],1942,4398,"PD-T7-1_WP_205975857.1,PD-T7-1_WP_205975857.1, 1, 2.3e-42, 0.977, 0.752 | PD-T7-5_WP_098786838.1,PD-T7-5_WP_098786838.1, 1, 1.4e-116, 0.977, 0.983","PD-T7-5_WP_098786838.1, PD-T7-5_WP_098786838.1, 1.4e-116, 0.977, 0.983 | PD-T7-1_WP_205975857.1, PD-T7-1_WP_205975857.1, 2.3e-42, 0.977, 0.752"
3,NZ_CP025084.1,Paris,WP_021015404.1,PDLC02979,AAA_15,AriA,9.7e-19,3.2e-18,0.919,0.96,3658314,3659795,+,AAA family ATPase [Serratia sp. ATCC 39006],3237,4398,"PDLC02979,AAA_15, 1, 3.2e-18, 0.919, 0.96 | PDLC02980,AAA_21, 1, 5.6e-16, 0.888, 0.977","PDLC02979, AAA_15, 3.2e-18, 0.919, 0.96 | PDLC02980, AAA_21, 5.6e-16, 0.888, 0.977"
3,NZ_CP025084.1,Paris,WP_021015403.1,PDLC02983,DUF4435,AriB,4.1e-19,5.7e-19,0.746,0.936,3659795,3660649,+,DUF4435 domain-containing protein [Serratia sp. ATCC 39006],3238,4398,"PDLC02983,DUF4435, 1, 5.7e-19, 0.746, 0.936","PDLC02983, DUF4435, 5.7e-19, 0.746, 0.936"
2,NZ_CP025084.1,Mokosh_TypeII,WP_021014804.1,Mokosh_TypeII__MkoC,Mokosh_TypeII__MkoC,MkoC,2.2999999999999996e-62,4.8999999999999995e-62,0.664,0.632,4364059,4367682,-,hypothetical protein [Serratia sp. ATCC 39006],3836,4398,"Mokosh_TypeII__MkoC,Mokosh_TypeII__MkoC, 1, 4.9e-62, 0.664, 0.632","Mokosh_TypeII__MkoC, Mokosh_TypeII__MkoC, 4.9e-62, 0.664, 0.632"
6,NZ_CP025084.1,SoFic,pseudo_subWP_004241487.1,SoFic__SoFic,SoFic__SoFic,SoFic,2.1999999999999997e-47,2.9999999999999997e-47,0.803,0.817,4444233,4445231,-,Fic family protein [Morganella morganii],3917,4398,"SoFic__SoFic,SoFic__SoFic, 1, 3e-47, 0.803, 0.817","SoFic__SoFic, SoFic__SoFic, 3e-47, 0.803, 0.817"
3,NZ_CP025084.1,PDC-S11,WP_021014227.1,PDLC04913,PDC-S11_WP_158522352.1,PDC-S11,1.0999999999999996e-175,1.2999999999999994e-175,0.957,0.992,24870,26057,+,DUF4268 domain-containing protein [Serratia sp. ATCC 39006],23,4398,"PDLC04909,PDC-S11_WP_104289981.1, 1, 6.2e-61, 0.901, 0.945 | PDLC04910,PDC-S11_WP_052717175.1, 1, 1.3e-57, 0.562, 0.599 | PDLC04911,PDC-S11_WP_167956302.1, 1, 2.5e-05, 0.228, 0.283 | PDLC04911,PDC-S11_WP_167956302.1, 2, 1.7e-28, 0.387, 0.481 | PDLC04912,PDC-S11_WP_055175232.1, 1, 0.0042, 0.228, 0.288 | PDLC04912,PDC-S11_WP_055175232.1, 2, 4.6e-25, 0.544, 0.668 | PDLC04913,PDC-S11_WP_158522352.1, 1, 1.3e-175, 0.957, 0.992 | PDLC04914,PDC-S11_WP_033147849.1, 1, 1e-06, 0.223, 0.271 | PDLC04914,PDC-S11_WP_033147849.1, 2, 1.6e-34, 0.4, 0.513 | PDLC04915,PDC-S11_WP_099259587.1, 1, 4.7e-53, 0.648, 0.652 | PDLC04916,PDC-S11_WP_098770551.1, 1, 4.7e-29, 0.529, 0.536","PDLC04913, PDC-S11_WP_158522352.1, 1.3e-175, 0.957, 0.992 | PDLC04909, PDC-S11_WP_104289981.1, 6.2e-61, 0.901, 0.945 | PDLC04910, PDC-S11_WP_052717175.1, 1.3e-57, 0.562, 0.599 | PDLC04915, PDC-S11_WP_099259587.1, 4.7e-53, 0.648, 0.652 | PDLC04914, PDC-S11_WP_033147849.1, 1.6e-34, 0.4, 0.513"
2,NZ_CP025084.1,PDC-S08,WP_021014224.1,PDLC04900,PDC-S08_WP_202707215.1,PDC-S08,4.3999999999999986e-133,5.099999999999998e-133,0.981,0.935,31798,32757,+,5'-nucleotidase [Serratia sp. ATCC 39006],26,4398,"PDLC04900,PDC-S08_WP_202707215.1, 1, 5.1e-133, 0.981, 0.935","PDLC04900, PDC-S08_WP_202707215.1, 5.1e-133, 0.981, 0.935"
1,NZ_CP025084.1,PDC-S07,WP_021017122.1,PDLC04899,PDC-S07_WP_110056698.1,PDC-S07,1.2e-36,1.3e-36,0.962,0.926,1345326,1345721,+,8-oxo-dGTP diphosphatase MutT [Serratia sp. ATCC 39006],1185,4398,"PDLC04899,PDC-S07_WP_110056698.1, 1, 1.3e-36, 0.962, 0.926","PDLC04899, PDC-S07_WP_110056698.1, 1.3e-36, 0.962, 0.926"
